magic
tech scmos
timestamp 1629535326
<< ntransistor >>
rect -48 -22 -46 -12
rect -30 -22 -28 -12
rect -12 -22 -10 -12
rect 6 -22 8 -12
<< ptransistor >>
rect -54 30 -34 32
rect -48 0 -46 20
rect -30 0 -28 20
rect -12 0 -10 20
rect 6 0 8 20
<< ndiffusion >>
rect -49 -22 -48 -12
rect -46 -22 -45 -12
rect -31 -22 -30 -12
rect -28 -22 -27 -12
rect -13 -22 -12 -12
rect -10 -22 -9 -12
rect 5 -22 6 -12
rect 8 -22 9 -12
<< pdiffusion >>
rect -54 32 -34 33
rect -54 29 -34 30
rect -49 0 -48 20
rect -46 0 -45 20
rect -31 0 -30 20
rect -28 0 -27 20
rect -13 0 -12 20
rect -10 0 -9 20
rect 5 0 6 20
rect 8 0 9 20
<< ndcontact >>
rect -54 -22 -49 -12
rect -45 -22 -40 -12
rect -36 -22 -31 -12
rect -27 -22 -22 -12
rect -18 -22 -13 -12
rect -9 -22 -4 -12
rect 0 -22 5 -12
rect 9 -22 14 -12
<< pdcontact >>
rect -54 33 -34 38
rect -54 24 -34 29
rect -54 0 -49 20
rect -45 0 -40 20
rect -36 0 -31 20
rect -27 0 -22 20
rect -18 0 -13 20
rect -9 0 -4 20
rect 0 0 5 20
rect 9 0 14 20
<< psubstratepcontact >>
rect -53 -38 -49 -34
rect -38 -38 -34 -34
rect -30 -38 -26 -34
rect -21 -38 -17 -34
rect -13 -38 -9 -34
rect -5 -38 -1 -34
rect 9 -38 13 -34
<< nsubstratencontact >>
rect -29 34 -25 38
rect -18 34 -14 38
rect -7 34 -3 38
rect 1 34 5 38
rect 10 34 14 38
<< polysilicon >>
rect -32 50 -14 52
rect -32 32 -30 50
rect -16 42 -14 50
rect -56 30 -54 32
rect -34 30 -30 32
rect -23 24 -21 42
rect -16 40 8 42
rect -58 21 -46 23
rect -48 20 -46 21
rect -30 22 -21 24
rect -13 22 -10 26
rect -30 20 -28 22
rect -12 20 -10 22
rect 6 20 8 40
rect -48 -2 -46 0
rect -30 -2 -28 0
rect -48 -8 -40 -5
rect -36 -8 -28 -5
rect -48 -12 -46 -8
rect -30 -12 -28 -8
rect -12 -12 -10 0
rect 6 -4 8 0
rect 0 -7 8 -4
rect 6 -12 8 -10
rect -48 -24 -46 -22
rect -30 -24 -28 -22
rect -12 -24 -10 -22
rect 6 -27 8 -22
rect -20 -30 8 -27
<< polycontact >>
rect -24 42 -20 46
rect -62 20 -58 24
rect -17 22 -13 26
rect -40 -8 -36 -4
rect -4 -8 0 -4
rect -24 -30 -20 -26
<< metal1 >>
rect -62 42 -24 46
rect -34 38 15 39
rect -34 34 -29 38
rect -25 34 -18 38
rect -14 34 -7 38
rect -3 34 1 38
rect 5 34 10 38
rect 14 34 15 38
rect -34 33 15 34
rect -45 20 -34 24
rect -18 26 -13 33
rect -18 22 -17 26
rect -18 20 -13 22
rect 0 20 5 33
rect -40 0 -36 20
rect -54 -4 -49 0
rect -54 -8 -40 -4
rect -54 -12 -49 -8
rect -27 -12 -22 0
rect -9 -12 -4 0
rect 9 -12 14 0
rect -45 -33 -40 -22
rect -36 -33 -31 -22
rect -26 -26 -22 -22
rect -26 -30 -24 -26
rect -17 -33 -13 -22
rect 0 -33 5 -22
rect -54 -34 14 -33
rect -54 -38 -53 -34
rect -49 -38 -38 -34
rect -34 -38 -30 -34
rect -26 -38 -21 -34
rect -17 -38 -13 -34
rect -9 -38 -5 -34
rect -1 -38 9 -34
rect 13 -38 14 -34
rect -54 -39 14 -38
<< labels >>
rlabel polycontact -60 22 -60 22 3 ninv
rlabel metal1 -60 44 -60 44 3 inv
rlabel metal1 -10 36 -10 36 1 vdd
rlabel metal1 3 -36 3 -36 1 vss
rlabel metal1 12 -6 12 -6 7 out
<< end >>
