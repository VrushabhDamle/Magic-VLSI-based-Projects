magic
tech scmos
timestamp 1621679198
<< ntransistor >>
rect 5 -22 7 -12
<< ptransistor >>
rect 5 0 7 20
<< ndiffusion >>
rect 4 -22 5 -12
rect 7 -22 9 -12
<< pdiffusion >>
rect 4 0 5 20
rect 7 0 9 20
<< ndcontact >>
rect 0 -22 4 -12
rect 9 -22 13 -12
<< pdcontact >>
rect 0 0 4 20
rect 9 0 13 20
<< psubstratepcontact >>
rect -3 -30 1 -26
rect 12 -30 16 -26
<< nsubstratencontact >>
rect -3 24 1 28
rect 12 24 16 28
<< polysilicon >>
rect 5 20 7 22
rect 5 -4 7 0
rect 3 -8 7 -4
rect 5 -12 7 -8
rect 5 -24 7 -22
<< polycontact >>
rect -1 -8 3 -4
<< metal1 >>
rect -4 28 17 29
rect -4 24 -3 28
rect 1 24 12 28
rect 16 24 17 28
rect -4 23 17 24
rect 0 20 4 23
rect 9 -12 13 0
rect 0 -25 4 -22
rect -4 -26 17 -25
rect -4 -30 -3 -26
rect 1 -30 12 -26
rect 16 -30 17 -26
rect -4 -31 17 -30
<< labels >>
rlabel metal1 3 25 3 25 5 vdd
rlabel metal1 3 -29 3 -29 1 gnd
rlabel metal1 11 -5 11 -5 1 Z
rlabel polycontact 1 -6 1 -6 3 A
<< end >>
