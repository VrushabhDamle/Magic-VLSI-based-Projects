magic
tech scmos
timestamp 1629385257
<< ntransistor >>
rect -12 -22 -10 -12
rect 6 -28 8 -18
rect 32 -28 34 -18
rect 50 -22 52 -12
<< ptransistor >>
rect 6 0 8 20
rect 32 0 34 20
<< ndiffusion >>
rect -13 -22 -12 -12
rect -10 -22 -9 -12
rect 5 -28 6 -18
rect 8 -28 9 -18
rect 31 -28 32 -18
rect 34 -28 35 -18
rect 49 -22 50 -12
rect 52 -22 53 -12
<< pdiffusion >>
rect 5 0 6 20
rect 8 0 9 20
rect 31 0 32 20
rect 34 0 35 20
<< ndcontact >>
rect -18 -22 -13 -12
rect -9 -22 -4 -12
rect 0 -28 5 -18
rect 9 -28 14 -18
rect 26 -28 31 -18
rect 35 -28 40 -18
rect 44 -22 49 -12
rect 53 -22 58 -12
<< pdcontact >>
rect 0 0 5 20
rect 9 0 14 20
rect 26 0 31 20
rect 35 0 40 20
<< psubstratepcontact >>
rect -16 -36 -12 -32
rect 1 -36 5 -32
rect 18 -36 22 -32
rect 35 -36 39 -32
rect 52 -36 56 -32
<< nsubstratencontact >>
rect 1 24 5 28
rect 18 24 22 28
rect 35 24 39 28
<< polysilicon >>
rect 6 20 8 22
rect 32 20 34 22
rect -12 -12 -10 -7
rect 6 -11 8 0
rect 32 -3 34 0
rect 22 -7 34 -3
rect 6 -15 18 -11
rect 6 -18 8 -15
rect 32 -18 34 -7
rect 50 -12 52 -7
rect -12 -24 -10 -22
rect 50 -24 52 -22
rect 6 -30 8 -28
rect 32 -30 34 -28
<< polycontact >>
rect -13 -7 -9 -3
rect 18 -7 22 -3
rect 49 -7 53 -3
rect 18 -15 22 -11
<< metal1 >>
rect -13 32 53 38
rect -27 -12 -21 20
rect -13 -3 -9 32
rect 0 28 40 29
rect 0 24 1 28
rect 5 24 18 28
rect 22 24 35 28
rect 39 24 40 28
rect 0 23 40 24
rect 9 20 14 23
rect 26 20 31 23
rect 0 -3 5 0
rect 0 -7 18 -3
rect 0 -12 5 -7
rect 35 -11 40 0
rect 49 -3 53 32
rect -27 -22 -18 -12
rect -4 -15 5 -12
rect 22 -12 40 -11
rect 61 -12 67 20
rect 22 -15 44 -12
rect 0 -18 5 -15
rect 35 -18 40 -15
rect -27 -28 -21 -22
rect 9 -31 14 -28
rect 58 -22 67 -12
rect 61 -28 67 -22
rect 26 -31 31 -28
rect -21 -32 61 -31
rect -21 -36 -16 -32
rect -12 -36 1 -32
rect 5 -36 18 -32
rect 22 -36 35 -32
rect 39 -36 52 -32
rect 56 -36 61 -32
rect -21 -37 61 -36
<< labels >>
rlabel metal1 10 26 10 26 1 vdd
rlabel metal1 10 -34 10 -34 1 gnd
rlabel metal1 20 35 20 35 5 wl
rlabel metal1 -24 -17 -24 -17 3 blz
rlabel metal1 64 -17 64 -17 7 bl
<< end >>
