magic
tech scmos
timestamp 1631598125
<< ntransistor >>
rect 5 -22 7 -12
<< ptransistor >>
rect 5 0 7 20
<< ndiffusion >>
rect 4 -22 5 -12
rect 7 -22 8 -12
<< pdiffusion >>
rect 4 0 5 20
rect 7 0 8 20
<< ndcontact >>
rect 0 -22 4 -12
rect 8 -22 12 -12
<< pdcontact >>
rect 0 0 4 20
rect 8 0 12 20
<< psubstratepcontact >>
rect -3 -30 1 -26
rect 11 -30 15 -26
<< nsubstratencontact >>
rect -3 24 1 28
rect 11 24 15 28
<< polysilicon >>
rect 5 20 7 22
rect 5 -4 7 0
rect 3 -8 7 -4
rect 5 -12 7 -8
rect 5 -24 7 -22
<< polycontact >>
rect -1 -8 3 -4
<< metal1 >>
rect -4 28 16 29
rect -4 24 -3 28
rect 1 24 11 28
rect 15 24 16 28
rect -4 23 16 24
rect 0 20 4 23
rect 8 -12 12 0
rect 0 -25 4 -22
rect -4 -26 16 -25
rect -4 -30 -3 -26
rect 1 -30 11 -26
rect 15 -30 16 -26
rect -4 -31 16 -30
<< labels >>
rlabel polycontact 1 -6 1 -6 3 A
rlabel metal1 10 -6 10 -6 1 Z
rlabel metal1 6 -28 6 -28 1 gnd
rlabel metal1 6 26 6 26 5 vdd
<< end >>
